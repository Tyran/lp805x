module lp805x_clk(rst,clki,sel,clko);

parameter CHOICES=4;

input 					rst;
input 					clki;
input [CHOICES-1:0] 	sel;

output					clko;





endmodule